library IEEE;
use IEEE.STD_LOGIC_1164.all;

package common is
	type carry_unit_t is (KOGGE_STONE, RIPPLE_CARRY);
end common;

package body common is
end common;
