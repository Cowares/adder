library IEEE;
use IEEE.STD_LOGIC_1164.all;

package common is
	type carry_unit_t is (BRENT_KUNG, HAN_CARLSON, KOGGE_STONE);
end common;

package body common is
end common;
