library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity KoggeStoneAdder is
	port (	
		P: in std_logic_vector;
		G: in std_logic_vector;
		cout: out std_logic
	);
end KoggeStoneAdder;

architecture Behavioral of KoggeStoneAdder is

begin


end Behavioral;
